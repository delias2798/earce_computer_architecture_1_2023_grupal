module memory #(parameter WIDTH=8)(
    input logic clk, reset, MemWriteM,
    input logic [WIDTH-1:0] ALUOutM, WriteData,
    output logic [WIDTH-1:0] ReadData
);

endmodule